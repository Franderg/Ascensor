`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:54:58 03/24/2017 
// Design Name: 
// Module Name:    manejo_entradas 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: maneja las entradas, convirtiendo lo que entra en un registro para
// poder ser usado por el resto del programa.
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module manejo_entradas(
    );


endmodule
